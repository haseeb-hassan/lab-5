module YourModule(input [3:0] num, input [2:0] set, output reg [6:0] w, output reg [7:0] y);
    always_comb begin
        case (num)
            4'b0000:  w = 7'b0000001;
            4'b0001:  w = 7'b1001111;
            4'b0010:  w = 7'b0010010;
            4'b0011:  w = 7'b0000110;
            4'b0100:  w = 7'b1001100;
            4'b0101:  w = 7'b0100100;
            4'b0110:  w = 7'b0100000;
            4'b0111:  w = 7'b0001111;
            4'b1000:  w = 7'b0000000;
            4'b1001:  w = 7'b0000100;
            4'b1010:  w = 7'b0001000;
            4'b1011:  w = 7'b1100000;
            4'b1100:  w = 7'b0110001;
            4'b1101:  w = 7'b1000010;
            4'b1110:  w = 7'b0110000;
            4'b1111:  w = 7'b0111000;
        endcase

        case (set)
            3'b000 : y = 8'b11111110;
            3'b001 : y = 8'b11111101;
            3'b010 : y = 8'b11111011;
            3'b011 : y = 8'b11110111;
            3'b100 : y = 8'b11101111;
            3'b101 : y = 8'b11011111;
            3'b110 : y = 8'b10111111;
            3'b111 : y = 8'b01111111;
            default : y = 8'b11111111;
        endcase 
    end
endmodule
